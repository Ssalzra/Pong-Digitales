LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

PACKAGE mtx_pkg IS 

TYPE Img_mtx IS ARRAY (0 TO 7) OF STD_LOGIC_VECTOR(15 DOWNTO 0);

END mtx_pkg;
